library ieee;
use ieee.numeric_bit.all;
use std.textio.all;

entity memoriaInstrucoes is
    generic (
        addressSize : natural := 8; -- Corrigido: removido espa�o em ": ="
        dataSize    : natural := 8; -- Corrigido: removido espa�o em ": ="
        datFileName : string  := "memInstr_conteudo.dat" -- Corrigido: removido espa�o em ": ="
    );
    port (
        addr : in  bit_vector(addressSize-1 downto 0);
        data : out bit_vector(dataSize-1 downto 0)
    );
end entity memoriaInstrucoes; -- Corrigido: nome deve bater com a declara��o

architecture mem_instru of memoriaInstrucoes is
    
    -- 1. Defini��o do Tipo deve vir ANTES da fun��o
    -- O tamanho agora � calculado com base no addressSize (2^N - 1)
    type mem_t is array (0 to (2**addressSize)-1) of bit_vector(dataSize-1 downto 0);

    -- 2. Fun��o de Inicializa��o
    impure function inicializa(nome_do_arquivo : in string) return mem_t is
        file     arquivo  : text open read_mode is nome_do_arquivo;
        variable linha    : line;
        variable temp_bv  : bit_vector(dataSize-1 downto 0);
        variable temp_mem : mem_t;
    begin
        -- Inicializa a mem�ria com zeros (boa pr�tica)
        temp_mem := (others => (others => '0'));
        
        for i in temp_mem'range loop
            if not endfile(arquivo) then
                readline(arquivo, linha);
                read(linha, temp_bv);
                temp_mem(i) := temp_bv;
            end if;
        end loop;
        return temp_mem;
    end function;

    -- 3. Declara��o dos Sinais
    signal mem      : mem_t := inicializa(datFileName);
    signal addr_int : natural; -- 'natural' � mais simples que integer range aqui

begin 
    -- 4. Convers�o correta usando numeric_bit
    -- bit_vector -> unsigned -> integer
    addr_int <= to_integer(unsigned(addr));
    
    -- Acesso � mem�ria
    data <= mem(addr_int);

end architecture mem_instru;